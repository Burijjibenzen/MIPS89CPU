`include "defines.vh"

module inst_rom( 
    input  wire               ce, 
    input  wire[`InstAddrBus] addr, 
    output reg [`InstBus]     inst 
); 
    // ����һ�����飬��С�� InstMemNum��Ԫ�ؿ���� InstBus 
    reg[`InstBus]  inst_mem[0 : `InstMemNum -1 ]; 
    
    // ʹ���ļ� inst_rom.data ��ʼ��ָ��洢�� 
    initial $readmemh ( "D:/TJU/ComputerSystem/MIPS89/inst_rom.data", inst_mem ); 
 
// ����λ�ź���Чʱ����������ĵ�ַ������ָ��洢�� ROM �ж�Ӧ��Ԫ�� 
always @ (*) begin 
    if (ce == `ChipDisable) begin 
        inst <= `ZeroWord; 
    end 
    else begin 
        inst <= inst_mem[addr[`InstMemNumLog2 + 1 : 2]]; 
        // �й�Ϊʲô���Բ��� PC ����ַΪ 0x00400000��
        // ��Ϊ��ַ����ֻȡ����ൽ�� 18 λ���Ǹ� ��4�� ����û��
        // ���ԸĲ��Ķ�û��Ӱ��
    end 
end 
 
endmodule