`timescale 1ns / 1ps

// main two part: 1.spi flash control 2. wb main bus
module flash_rom(
    // Wishbone ���߽ӿ�
    input wire wb_clk_i,        // Wishbone ʱ��
    input wire wb_rst_i,        // Wishbone ��λ
    input wire wb_cyc_i,        // Wishbone ����������Ч
    input wire wb_stb_i,        // Wishbone ѡͨ�ź�
    input wire wb_we_i,         // Wishbone дʹ��
    input wire [3:0] wb_sel_i,  // Wishbone �ֽ�ѡ��
    input wire [23:0] wb_adr_i, // Wishbone ��ַ
    input wire [31:0] wb_dat_i, // Wishbone д����
    output reg [31:0] wb_dat_o, // Wishbone ������
    output reg        wb_ack_o, // Wishbone Ӧ��

    input wire flash_continue, // Flash ���������ź�

    // SPI Flash �ӿ�
    output reg cs_n,   // Ƭѡ�źţ�����Ч
    input  sdi,        // SPI �������루�� Flash �� FPGA��
    output reg sdo,    // SPI ����������� FPGA �� Flash��
    output reg wp_n,   // д����������Ч
    output reg hld_n   // �����źţ�����Ч
    );


// ״̬��״̬����
parameter IDLE       = 5'b00000;
parameter START      = 5'b00010;
parameter INST_OUT   = 5'b00011;
parameter ADDR1_OUT  = 5'b00100;
parameter ADDR2_OUT  = 5'b00101;
parameter ADDR3_OUT  = 5'b00110;
parameter WRITE_DATA = 5'b00111;
parameter READ_DATA  = 5'b01000;
parameter READ_DATA1 = 5'b01001;
parameter READ_DATA2 = 5'b01010;
parameter READ_DATA3 = 5'b01011;
parameter READ_DATA4 = 5'b01100;
parameter READ_DATA5 = 5'b01101;
parameter WAITING    = 5'b10000;
parameter ENDING     = 5'b10001;


// ��ʼ��������
(* dont_touch = "true" *)reg[4:0] init_count;

// SPI ������ؼĴ���
(* dont_touch = "true" *)reg         sck;        // SPI ʱ��
(* dont_touch = "true" *)reg  [4:0]  state;      // ��ǰ״̬
reg  [4:0]  next_state;                         // ��һ��״̬

(* dont_touch = "true" *)reg  [7:0]   instruction;   // SPI ָ��
(* dont_touch = "true" *)reg  [7:0]   datain_shift;  // SPI ������λ�Ĵ���
(* dont_touch = "true" *)reg  [7:0]   datain;        // SPI ��������
(* dont_touch = "true" *)reg  [7:0]   dataout;       // SPI �������
(* dont_touch = "true" *)reg          sck_en;        // SPI ʱ��ʹ��
(* dont_touch = "true" *)reg  [2:0]   sck_en_d;      // SPI ʱ��ʹ���ӳ�
(* dont_touch = "true" *)reg [10:0]   read_count;    // ��������
reg  [2:0]  cs_n_d;                                 // Ƭѡ�ź��ӳ�

reg         temp;                                   // ��ʱ����
(* dont_touch = "true" *)reg  [3:0]  sdo_count;     // SPI �������
reg  [15:0] page_count;                             // ҳ����
reg  [7:0]  wait_count;                             // �ȴ�����
(* dont_touch = "true" *)reg  [23:0] addr;          // 24 λ��ַ
reg         wrh_rdl;                                // д/����־��1 Ϊд��0 Ϊ��
reg         addr_req;                               // ��ַ�����־
reg  [15:0] wr_cnt;                                 // д�ֽ���
reg  [15:0] rd_cnt;                                 // ���ֽ���
(* dont_touch = "true" *)reg [31:0] read_data;      // ����������


// ״̬����Wishbone �ӿ��� SPI Flash����
always @ (posedge wb_clk_i or posedge wb_rst_i) begin
    if(wb_rst_i) begin
        // �첽��λ�����йؼ��Ĵ�����ʼ��
        state      <= IDLE;        // ״̬���ص� IDLE ����״̬
        read_count <= 11'd0;       // ����������
        wb_ack_o   <= 1'b0;        // Wishbone Ӧ���ź�����
        init_count <= 5'd2;        // ��ʼ��������
    end
    else if(wb_cyc_i & wb_stb_i) begin
        // Wishbone ������Чʱ��״̬���л�����һ��״̬
        state <= next_state;
        // �����ǰ���� ENDING ״̬�һ�δӦ��
        if(state == ENDING && !wb_ack_o) begin
            if(init_count > 5'd0) begin
                // �ӳ�һ��ʱ���ص� IDLE����ֹ���߳�ͻ
                init_count <= init_count - 5'd1;
                state      <= IDLE;
            end
            else 
                wb_ack_o   <= 1'b1; // ���ո���Ӧ���ź�
        end
    end
    else begin
        // Wishbone ��Чʱ��״̬���ص� IDLE��Ӧ���ź�����
        state    <= IDLE;
        wb_ack_o <= 1'b0;
    end
end

// SPI �����ź�Ĭ��ֵ����
always @ (posedge wb_clk_i) begin
    // ÿ��ʱ�����ڶ���д�����ͱ����ź����ߣ���ʹ�ܣ�
    wp_n  <= 1'b1;
    hld_n <= 1'b1;
end


// ״̬�������̼���״̬�¼Ĵ�����ֵ
always @ (posedge wb_clk_i or posedge wb_rst_i) begin
	if(wb_rst_i) begin
		// �첽��λ������ SPI ��ؼĴ�����ʼ��
        next_state  <= IDLE;      // ��һ��״̬Ϊ IDLE
        sck_en      <= 1'b0;      // SPI ʱ�ӽ�ֹ
        cs_n_d[0]   <= 1'b1;      // Ƭѡ���ߣ���ѡ�У�
        dataout     <= 8'd0;      // SPI �����������
        sdo_count   <= 4'd0;      // SPI �����������
        sdo         <= 1'b0;      // SPI �������������
        datain      <= 8'd0;      // SPI ������������
        addr        <=24'd0;      // ��ַ����
        datain_shift<=8'd0;       // ������λ�Ĵ�������
        temp        <= 1'b0;      // ��ʱ��������
        page_count  <= 16'd0;     // ҳ��������
        wait_count  <= 8'd0;      // �ȴ���������
        read_data   <=32'd0;      // �����ݼĴ�������
        
	end
	else begin
		case(state)
		// ����״̬���ȴ� flash_continue �ź����ߺ���� START
		IDLE: 
		begin
            wait_count <= 8'd0; // �ȴ���������
            if(flash_continue==1'd1)
                next_state<=START; // ��⵽ flash_continue �źţ�׼������ SPI
            // ���򱣳��� IDLE
        end
		
		START:
		// ����״̬��׼�� SPI ͨ�ţ����� CS�����ص�ַ
		begin
            addr       <= wb_adr_i;      // ���� Wishbone ����� 24 λ��ַ
            sck_en     <= 1'b1;      // ʹ�� SPI ʱ��
            cs_n_d[0]  <= 1'b0;  // ����Ƭѡ��ѡ�� Flash
            next_state <= INST_OUT; // ����ָ���״̬
            read_count <= read_count + 11'd1; // ������ +1
        end

		// ָ���״̬���� 8 λ SPI ָ����λ�Ƴ�
        INST_OUT:
        begin
            // sdo_count == 1 ʱ������ָ���λ�Ĵ���
            if(sdo_count == 4'd1) begin
                {sdo, dataout[6:0]} <= instruction;
            end
            // �����������ڣ���λ���
            else if(sdo_count[0]) begin
                {sdo, dataout[6:0]} <= {dataout[6:0], 1'b0};
            end

            // ������ 16 ��ʱ�ӣ�8 λ���� +8 ����ʱ�ӣ�������
            if(sdo_count != 4'd15) begin
                sdo_count <= sdo_count + 4'd1;
            end
            else begin
                sdo_count  <= 4'd0;
                // �ж��Ƿ���Ҫ����ַ������ֱ�ӽ������ݽ׶�
                next_state <= (addr_req) ?  ADDR1_OUT : ((wrh_rdl) ? ((wr_cnt==16'd0) ? ENDING : WRITE_DATA) : ((rd_cnt==16'd0) ? ENDING : READ_DATA1));
            end
        end

		// ���͵�ַ�� 8 λ
        ADDR1_OUT:
        begin
            if(sdo_count == 4'd1) begin
                {sdo, dataout[6:0]} <= addr[23:16];
            end
            else if(sdo_count[0]) begin
                {sdo, dataout[6:0]} <= {dataout[6:0],1'b0};
            end

            if(sdo_count != 4'd15) begin
                sdo_count <= sdo_count + 4'd1;
            end
            else begin
                sdo_count  <= 4'd0;
                next_state <= ADDR2_OUT; // ������ 8 λ��ַ����
            end
        end

		// ���͵�ַ�� 8 λ
        ADDR2_OUT:
        begin
            if(sdo_count == 4'd1) begin
                {sdo, dataout[6:0]} <= addr[15:8];
            end
            else if(sdo_count[0]) begin
                {sdo, dataout[6:0]} <= {dataout[6:0], 1'b0};
            end

            if(sdo_count != 4'd15) begin
                sdo_count <= sdo_count + 4'd1;
            end
            else begin
                sdo_count  <= 4'd0;
                next_state <= ADDR3_OUT; // ����� 8 λ��ַ����
            end
        end

		// ���͵�ַ�� 8 λ
        ADDR3_OUT:
        begin
            if(sdo_count == 4'd1) begin
                {sdo, dataout[6:0]} <= addr[7:0];
            end
            else if(sdo_count[0]) begin
                {sdo, dataout[6:0]} <= {dataout[6:0], 1'b0};
            end

            if(sdo_count != 4'd15) begin
                sdo_count <= sdo_count + 4'd1;
            end
            else begin
                sdo_count  <= 4'd0;
                // �ж���д���Ƕ�
                next_state <= (wrh_rdl) ? ((wr_cnt==16'd0) ? ENDING : WRITE_DATA) : ((rd_cnt==16'd0) ? ENDING : READ_DATA1);
                page_count <= 16'd0; // ҳ��������
            end
        end

		// д����״̬������Ϊ�������� 0x5A��
        WRITE_DATA:
        begin
            if(sdo_count == 4'd1) begin
                {sdo, dataout[6:0]} <= 8'h5A;
            end
            else if(sdo_count[0]) begin
                {sdo, dataout[6:0]} <= {dataout[6:0], 1'b0};
            end

            if(sdo_count != 4'd15) begin
                sdo_count <= sdo_count + 4'd1;
            end
            else begin
                page_count <= page_count + 16'd1;
                sdo_count  <= 4'd0;
                // �ж��Ƿ�д����������
                next_state <= (page_count < (wr_cnt - 16'd1)) ? WRITE_DATA : ENDING;
            end
        end

		// �����ݵ� 1 �ֽڣ������ֽڣ�����λ����
        READ_DATA1:
        begin
            // ż��������λ���� sdi
            if(~sdo_count[0]) begin
                datain_shift <= {datain_shift[6:0], sdi};
            end
            // sdo_count == 1 ʱ������� 1 �ֽ�
            if(sdo_count == 4'd1) begin
                datain <= {datain_shift, sdi};
            end

            if(sdo_count != 4'd15) begin
                sdo_count <= sdo_count + 4'd1;
            end
            else begin
                page_count <= page_count + 16'd1;
                sdo_count  <= 4'd0;
                next_state <= READ_DATA2; // ����� 2 �ֽڽ���
            end
        end

        READ_DATA2: // ֻ�����µ� 2 �����������Ե�ǰ���ڴ���� SPI �ֽ����ģ����� 6 �������ǡ��¾ɡ���
        begin
            if(~sdo_count[0]) begin
                datain_shift <= {datain_shift[6:0], sdi};
            end
            if(sdo_count == 4'd1) begin
                read_data[31:24] <= {datain_shift, sdi};
                datain<= {datain_shift, sdi};
            end

            if(sdo_count != 4'd15) begin
                sdo_count <= sdo_count + 4'd1;
            end
            else begin
                page_count <= page_count + 16'd1;
                sdo_count  <= 4'd0;
                next_state <= READ_DATA3; // ����� 3 �ֽڽ���
            end
        end

		// �����ݵ� 3 �ֽڣ����� read_data[23:16]
        READ_DATA3:
        begin
            if(~sdo_count[0]) begin
                datain_shift <= {datain_shift[6:0],sdi};
            end
            if(sdo_count == 4'd1) begin
                read_data[23:16] <= {datain_shift, sdi};
                datain<= {datain_shift, sdi};
            end

            if(sdo_count != 4'd15) begin
                sdo_count <= sdo_count + 4'd1;
            end
            else begin
                page_count <= page_count + 16'd1;
                sdo_count  <= 4'd0;
                next_state <=READ_DATA4; // ����� 4 �ֽڽ���
            end
        end

		// �����ݵ� 4 �ֽڣ����� read_data[15:8]
        READ_DATA4:
        begin
            if(~sdo_count[0]) begin
                datain_shift <= {datain_shift[6:0],sdi};
            end
            if(sdo_count == 4'd1) begin
                read_data[15:8] <= {datain_shift, sdi};
                datain<= {datain_shift, sdi};
            end

            if(sdo_count != 4'd15) begin
                sdo_count <= sdo_count + 4'd1;
            end
            else begin
                page_count <= page_count + 16'd1;
                sdo_count  <= 4'd0;
                next_state <=READ_DATA5; // ����� 5 �ֽڽ���
            end
        end

		// �����ݵ� 5 �ֽڣ����� read_data[7:0]
        READ_DATA5:
        begin
            if(~sdo_count[0]) begin
                datain_shift <= {datain_shift[6:0],sdi};
            end
            if(sdo_count == 4'd1) begin
                read_data[7:0] <= {datain_shift, sdi};
                datain<= {datain_shift, sdi};
            end

            if(sdo_count != 4'd15) begin
                sdo_count <= sdo_count + 4'd1;
            end
            else begin
                page_count <= page_count + 16'd1;
                sdo_count  <= 4'd0;
                next_state <=WAITING; // ���ݽ�����ϣ�����ȴ�
            end
        end

		// �ȴ�״̬���ر� SCK �� CS��׼������
        WAITING:
        begin
            sck_en <= 1'b0;      // ��ֹ SPI ʱ��
            cs_n_d[0] <= 1'b1;   // ����Ƭѡ���ͷ� Flash
            sdo_count <= 4'd0;   // �����������
            next_state<=ENDING;  // �������״̬
        end

		// ����״̬���ȴ� Wishbone Ӧ��
        ENDING:
        begin
            // �գ��ȴ��ⲿ always �鴦��Ӧ���ź�
        end
		endcase
	end
end

// SCK ������������ SPI ʱ���ź�
always @ (posedge wb_clk_i) begin
    // sck_en_d �� sck_en �Ĵ����ӳ٣�����ͬ���ͱ��ؼ��
    sck_en_d <= {sck_en_d[1:0], sck_en};
end

always @ (posedge wb_clk_i or posedge wb_rst_i) begin
    if(wb_rst_i) begin
        sck <= 1'b0; // ��λʱ SPI ʱ������
    end
    // sck_en_d[2] & sck_en Ϊ��ʱ����ת sck��ʵ�� SPI ʱ��
    else if(sck_en_d[2] & sck_en) begin
        sck <= ~sck;
    end
    else begin
        sck <= 1'b0; // ����������ֵ͵�ƽ
    end
end

// Ƭѡ�ź��ӳٴ�����֤ SPI ʱ���ȶ�
always @ (posedge wb_clk_i or posedge wb_rst_i) begin
    if(wb_rst_i) begin
        {cs_n, cs_n_d[2:1]} <= 3'h7; // ��λʱƬѡ���ߣ���ѡ�У�
    end
    else begin
        {cs_n, cs_n_d[2:1]} <= cs_n_d; // Ƭѡ�ź���λ���ӳ����
    end
end

// STARTUPE2 ԭ����ڽ��û�ʱ�ӣ�sck������� SPI Flash �� SCK ����
STARTUPE2
#(
.PROG_USR("FALSE"),
.SIM_CCLK_FREQ(10.0)
)
STARTUPE2_inst
(
  .CFGCLK     (),           // δ��
  .CFGMCLK    (),           // δ��
  .EOS        (),           // δ��
  .PREQ       (),           // δ��
  .CLK        (1'b0),       // δ��
  .GSR        (1'b0),       // δ��
  .GTS        (1'b0),       // δ��
  .KEYCLEARB  (1'b0),       // δ��
  .PACK       (1'b0),       // δ��
  .USRCCLKO   (sck),        // �û� SPI ʱ�����
  .USRCCLKTS  (1'b0),       // 0 ʹ�� CCLK ���
  .USRDONEO   (1'b1),       // 1
  .USRDONETS  (1'b1)        // 1
);

// ָ��������������ã�����Ϊ�̶���ָ�
always @ (posedge wb_clk_i) begin
    instruction <= 8'h03;    // ��ָ�0x03��
    wrh_rdl     <= 1'b0;     // ������
    addr_req    <= 1'b1;     // ��Ҫ���͵�ַ
    wr_cnt      <= 16'd0;    // д�ֽ���Ϊ0
    rd_cnt      <= 16'd4;    // ��4�ֽ�
end

// Wishbone ���������
always @ (posedge wb_clk_i) begin
    wb_dat_o <= read_data;   // ����ȡ������������� Wishbone ����
end
 
endmodule