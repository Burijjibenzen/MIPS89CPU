module wishbone_bus_if(
    input  wire        clk,    
    input  wire        rst, 
    
    // ���� ctrl ģ�� 
    input  wire[5:0]              stall_i, 
    input  wire                   flush_i,     // �����쳣����Ҫ�����ˮ��
    
    // CPU ��Ľӿ� 
    input  wire                   cpu_ce_i,    // ���Դ������ķ��������ź�
    input  wire[`RegBus]          cpu_data_i,  // ���Դ�����������
    input  wire[`RegBus]          cpu_addr_i, 
    input  wire                   cpu_we_i, 
    input  wire[3:0]              cpu_sel_i, 
    output reg[`RegBus]           cpu_data_o,  // ����������������� 
    
    // Wishbone ��Ľӿ� 
    input  wire[`RegBus]          wishbone_data_i,  // Wishbone �������������
    input  wire                   wishbone_ack_i, 
    output reg[`RegBus]           wishbone_addr_o, 
    output reg[`RegBus]           wishbone_data_o, 
    output reg                    wishbone_we_o, 
    output reg[3:0]               wishbone_sel_o, 
    output reg                    wishbone_stb_o,   // Wishbone ����ѡͨ�ź� 
    output reg                    wishbone_cyc_o,   // Wishbone ���������ź� 
    
    output reg                    stallreq  
);

    reg[1:0]     wishbone_state;   // ���� Wishbone ���߽ӿ�ģ���״̬ 
    reg[`RegBus] rd_buf;           // �Ĵ�ͨ�� Wishbone ���߷��ʵ������� 

/**************************************************************** 
***********          ��һ�Σ�����״̬ת����ʱ���·         ********* 
*****************************************************************/ 

always @ (posedge clk) begin 
    if(rst == `RstEnable) begin 
        wishbone_state  <= `WB_IDLE;         // ���� WB_IDLE ״̬ 
        wishbone_addr_o <= `ZeroWord; 
        wishbone_data_o <= `ZeroWord; 
        wishbone_we_o   <= `WriteDisable; 
        wishbone_sel_o  <= 4'b0000; 
        wishbone_stb_o  <= 1'b0;
        wishbone_cyc_o  <= 1'b0; 
        rd_buf          <= `ZeroWord; 
    end 
    else begin 
        case (wishbone_state) 
            `WB_IDLE: begin              // WB_IDLE ״̬ 
                if((cpu_ce_i == 1'b1) && (flush_i == `False_v)) begin 
                    wishbone_stb_o  <= 1'b1; 
                    wishbone_cyc_o  <= 1'b1; 
                    wishbone_addr_o <= cpu_addr_i; 
                    wishbone_data_o <= cpu_data_i; 
                    wishbone_we_o   <= cpu_we_i; 
                    wishbone_sel_o  <= cpu_sel_i; 
                    wishbone_state  <= `WB_BUSY;    // ���� WB_BUSY ״̬ 
                    rd_buf          <= `ZeroWord; 
                end 
            end 
            `WB_BUSY: begin              // WB_BUSY ״̬ 
                if(wishbone_ack_i == 1'b1) begin    // �յ� Wishbone ���ߵ���Ӧ
                    wishbone_stb_o  <= 1'b0; 
                    wishbone_cyc_o  <= 1'b0; 
                    wishbone_addr_o <= `ZeroWord; 
                    wishbone_data_o <= `ZeroWord; 
                    wishbone_we_o   <= `WriteDisable; 
                    wishbone_sel_o  <= 4'b0000; 
                    wishbone_state  <= `WB_IDLE;     // ���� WB_IDLE ״̬ 
                    if(cpu_we_i == `WriteDisable) begin  // ��ʾ������
                        rd_buf <= wishbone_data_i;       // �����������ݱ��浽���� rd_buf ��
                    end 
                    if(stall_i != 6'b000000) begin   // ��ˮ���в�����ͣ��
                    // ���� WB_WAIT_FOR_STALL ״̬ 
                        wishbone_state <= `WB_WAIT_FOR_STALL; 
                    end      
                end 
                else if(flush_i == `True_v) begin    // �ڻ�û���յ� Wishbone ���ߵ���Ӧʱ���������쳣
                    wishbone_stb_o  <= 1'b0; 
                    wishbone_cyc_o  <= 1'b0; 
                    wishbone_addr_o <= `ZeroWord; 
                    wishbone_data_o <= `ZeroWord; 
                    wishbone_we_o   <= `WriteDisable; 
                    wishbone_sel_o  <=  4'b0000; 
                    wishbone_state  <= `WB_IDLE;     // ���� WB_IDLE ״̬ 
                    rd_buf          <= `ZeroWord; 
                end 
            end 
            `WB_WAIT_FOR_STALL:  begin    // WB_WAIT_FOR_STALL ״̬ 
                if(stall_i == 6'b000000) begin   // ��ˮ����ͣ����
                    wishbone_state <= `WB_IDLE;   // ���� WB_IDLE ״̬ 
                end 
            end 
            default: begin 
            end  
        endcase 
    end    // if 
end      // always

/**************************************************************** 
***********      �ڶ��Σ����������ӿ��źŸ�ֵ����ϵ�·      ********* 
*****************************************************************/ 
always @ (*) begin 
    if(rst == `RstEnable) begin 
        stallreq   <= `NoStop; 
        cpu_data_o <= `ZeroWord; 
    end 
    else begin 
        stallreq   <= `NoStop; 
        case (wishbone_state) 
            `WB_IDLE: begin         // WB_IDLE ״̬ 
                if((cpu_ce_i == 1'b1) && (flush_i == `False_v)) begin  // ������Ҫ�������ߣ���û�д�����ˮ�����������
                    stallreq   <= `Stop;      // ��ͣ��ˮ���Եȴ��˴� Wishbone ���߷��ʽ���
                    cpu_data_o <= `ZeroWord; 
                end 
            end 
            `WB_BUSY: begin         // WB_BUSY ״̬ 
                if(wishbone_ack_i == 1'b1) begin  // �յ� Wishbone ���ߵ���Ӧ
                    stallreq <= `NoStop;          // ��ˮ�߿��Լ���
                    if(wishbone_we_o == `WriteDisable) begin  // ������
                        cpu_data_o <= wishbone_data_i;  // �� Wishbone ���߶��������ݴ��ݸ�������
                    end 
                    else begin 
                        cpu_data_o <= `ZeroWord; 
                    end 
                end 
                else begin                        // û���յ� Wishbone ���ߵ���Ӧ
                    stallreq   <= `Stop; 
                    cpu_data_o <= `ZeroWord;      // �˴η��ʻ�û�н�������ˮ��Ҫ������ͣ
                end 
            end 
            `WB_WAIT_FOR_STALL: begin  // WB_WAIT_FOR_STALL ״̬ 
                stallreq   <= `NoStop;            // Wishbone ���߷����Ѿ�����
                cpu_data_o <= rd_buf; 
            end 
            default: begin 
            end  
        endcase 
    end 
end

endmodule
