module mem(
    input wire              rst, 
    
    // ����ִ�н׶ε���Ϣ  
    input wire[`RegAddrBus] wd_i, 
    input wire              wreg_i, 
    input wire[`RegBus]     wdata_i, 
    input wire[`RegBus]     hi_i, 
    input wire[`RegBus]     lo_i, 
    input wire              whilo_i,
    
    input wire[`AluOpBus]   aluop_i,     // �ô�׶ε�ָ��Ҫ���е������������
    input wire[`RegBus]     mem_addr_i,  // �ô�׶εļ��ء��洢ָ���Ӧ�Ĵ洢����ַ
    input wire[`RegBus]     reg2_i,      // �ô�׶εĴ洢ָ��Ҫ�洢�����ݣ����� lwl��lwr ָ��Ҫд���Ŀ�ļĴ�����ԭʼֵ
    
    // �����ⲿ���ݴ洢�� RAM ����Ϣ�������ݴ洢����ȡ������
    input wire[`RegBus]     mem_data_i,  // �洢���� 32 λ��ַ��ÿ����ַ�� 1 �ֽ�
    
    input wire              LLbit_i,           // LLbit ģ������� LLbit �Ĵ�����ֵ
    input wire              wb_LLbit_we_i,     // ��д�׶ε�ָ���Ƿ�Ҫд LLbit �Ĵ��� 
    input wire              wb_LLbit_value_i,  // ��д�׶�Ҫд�� LLbit �Ĵ�����ֵ
    
    input wire              cp0_reg_we_i, 
    input wire[4:0]         cp0_reg_write_addr_i, 
    input wire[`RegBus]     cp0_reg_data_i,
    
    // ����ִ�н׶�
    input wire[31:0]        excepttype_i, 
    input wire              is_in_delayslot_i, 
    input wire[`RegBus]     current_inst_address_i,
    
    // ���� CP0 ģ��
    input wire[`RegBus]     cp0_status_i, 
    input wire[`RegBus]     cp0_cause_i, 
    input wire[`RegBus]     cp0_epc_i,
    
    // ���Ի�д�׶Σ��ǻ�д�׶ε�ָ��� CP0 �мĴ�����д��Ϣ�� 
    // �������������� 
    input wire              wb_cp0_reg_we, 
    input wire[4:0]         wb_cp0_reg_write_addr, 
    input wire[`RegBus]     wb_cp0_reg_data,
    
    // �ô�׶εĽ�� 
    output reg[`RegAddrBus] wd_o, 
    output reg              wreg_o, 
    output reg[`RegBus]     wdata_o,
    output reg[`RegBus]     hi_o, 
    output reg[`RegBus]     lo_o, 
    output reg              whilo_o,
    
    // �͵��ⲿ���ݴ洢��RAM����Ϣ
    output reg[`RegBus]     mem_addr_o,  // Ҫ���ʵ����ݴ洢���ĵ�ַ
    output wire             mem_we_o,    // �Ƿ���д������Ϊ 1 ��ʾ��д����
    output reg[3:0]         mem_sel_o,   // �ֽ�ѡ���ź�
    output reg[`RegBus]     mem_data_o,  // Ҫд�����ݴ洢��������
    output reg              mem_ce_o,    // ���ݴ洢��ʹ���ź�
    output reg              LLbit_we_o,     // �ô�׶ε�ָ���Ƿ�Ҫд LLbit �Ĵ���
    output reg              LLbit_value_o,  // �ô�׶ε�ָ��Ҫд�� LLbit �Ĵ�����ֵ
    
    output reg              cp0_reg_we_o, 
    output reg[4:0]         cp0_reg_write_addr_o, 
    output reg[`RegBus]     cp0_reg_data_o,
    
    output reg[31:0]        excepttype_o,       // ���յ��쳣����
    output wire[`RegBus]    cp0_epc_o,          // CP0 �� EPC �Ĵ���������ֵ
    output wire             is_in_delayslot_o,  // �ô�׶ε�ָ���Ƿ����ӳٲ�ָ��

    output wire[`RegBus]    current_inst_address_o // �ô�׶�ָ��ĵ�ַ
);

    reg               LLbit;      // ���� LLbit �Ĵ���������ֵ

    reg[`RegBus]      cp0_status;   // �������� CP0 �� Status �Ĵ���������ֵ 
    reg[`RegBus]      cp0_cause;    // �������� CP0 �� Cause �Ĵ���������ֵ 
    reg[`RegBus]      cp0_epc;      // �������� CP0 �� EPC �Ĵ���������ֵ 

    wire[`RegBus]     zero32; 
    reg               mem_we; 
 
    assign zero32   = `ZeroWord;
    
    // is_in_delayslot_o ��ʾ�ô�׶ε�ָ���Ƿ����ӳٲ�ָ�� 
    assign is_in_delayslot_o = is_in_delayslot_i;
    
    // current_inst_address_o �Ƿô�׶�ָ��ĵ�ַ 
    assign current_inst_address_o = current_inst_address_i;
    
  // ��ȡ LLbit �Ĵ���������ֵ�������д�׶ε�ָ��Ҫд LLbit����ô��д�׶�Ҫд��� 
  // ֵ���� LLbit �Ĵ���������ֵ����֮��LLbit ģ�������ֵ LLbit_i ������ֵ 
always @ (*) begin 
    if(rst == `RstEnable) begin 
        LLbit <= 1'b0; 
    end 
    else begin 
        if(wb_LLbit_we_i == 1'b1) begin 
            LLbit <= wb_LLbit_value_i;     // ��д�׶ε�ָ��Ҫд LLbit 
        end 
        else begin 
            LLbit <= LLbit_i; 
        end 
    end 
end

always @ (*) begin 
    if(rst == `RstEnable) begin 
        wd_o    <= `NOPRegAddr; 
        wreg_o  <= `WriteDisable; 
        wdata_o <= `ZeroWord; 
        hi_o    <= `ZeroWord; 
        lo_o    <= `ZeroWord; 
        whilo_o <= `WriteDisable;
        mem_addr_o <= `ZeroWord; 
        mem_we     <= `WriteDisable; 
        mem_sel_o  <= 4'b0000; 
        mem_data_o <= `ZeroWord; 
        mem_ce_o   <= `ChipDisable;
        LLbit_we_o    <= 1'b0; 
        LLbit_value_o <= 1'b0;
        cp0_reg_we_o         <= `WriteDisable; 
        cp0_reg_write_addr_o <= 5'b00000; 
        cp0_reg_data_o       <= `ZeroWord;
    end 
    else begin 
        wd_o    <= wd_i; 
        wreg_o  <= wreg_i; 
        wdata_o <= wdata_i; 
        hi_o    <= hi_i; 
        lo_o    <= lo_i; 
        whilo_o <= whilo_i;
        LLbit_we_o    <= 1'b0; 
        LLbit_value_o <= 1'b0;
        mem_we     <= `WriteDisable; 
        mem_addr_o <= `ZeroWord; 
        mem_sel_o  <= 4'b1111; 
        mem_ce_o   <= `ChipDisable;
        // ���� CP0 �мĴ�����д��Ϣ���ݵ���ˮ����һ�� 
        cp0_reg_we_o         <= cp0_reg_we_i; 
        cp0_reg_write_addr_o <= cp0_reg_write_addr_i; 
        cp0_reg_data_o       <= cp0_reg_data_i;
        
        case (aluop_i)
            `EXE_LB_OP: begin                  // lb ָ�� 
                mem_addr_o <= mem_addr_i; 
                mem_we     <= `WriteDisable; 
                mem_ce_o   <= `ChipEnable; 
                case (mem_addr_i[1:0]) 
                    2'b00: begin 
                        wdata_o   <= {{24{mem_data_i[31]}}, mem_data_i[31:24]};  // �͵�ַ
                        mem_sel_o <= 4'b1000; // ָ���� ��������ֵĵ�һ���ֽ�
                    end 
                    2'b01: begin 
                        wdata_o   <= {{24{mem_data_i[23]}}, mem_data_i[23:16]}; 
                        mem_sel_o <= 4'b0100; // ָ���� ��������ֵĵڶ����ֽ�
                    end 
                    2'b10: begin 
                        wdata_o   <= {{24{mem_data_i[15]}}, mem_data_i[15:8]}; 
                        mem_sel_o <= 4'b0010; 
                    end 
                    2'b11: begin 
                        wdata_o   <= {{24{mem_data_i[7]}}, mem_data_i[7:0]};    // �ߵ�ַ
                        mem_sel_o <= 4'b0001; 
                    end 
                    default: begin 
                        wdata_o   <= `ZeroWord; 
                    end 
                endcase 
            end
            `EXE_LBU_OP: begin            // lbu ָ�� 
                mem_addr_o <= mem_addr_i; 
                mem_we     <= `WriteDisable; 
                mem_ce_o   <= `ChipEnable; 
                case (mem_addr_i[1:0]) 
                    2'b00: begin 
                        wdata_o   <= {{24{1'b0}}, mem_data_i[31:24]}; 
                        mem_sel_o <= 4'b1000; 
                    end 
                    2'b01: begin 
                        wdata_o   <= {{24{1'b0}}, mem_data_i[23:16]}; 
                        mem_sel_o <= 4'b0100; 
                    end
                    2'b10: begin 
                        wdata_o   <= {{24{1'b0}}, mem_data_i[15:8]}; 
                        mem_sel_o <= 4'b0010; 
                    end 
                    2'b11: begin 
                        wdata_o   <= {{24{1'b0}}, mem_data_i[7:0]}; 
                        mem_sel_o <= 4'b0001; 
                    end 
                    default: begin 
                        wdata_o   <= `ZeroWord; 
                    end 
                endcase 
            end
            `EXE_LH_OP: begin                  // lh ָ�� 
                mem_addr_o <= mem_addr_i; 
                mem_we     <= `WriteDisable; 
                mem_ce_o   <= `ChipEnable; 
                case (mem_addr_i[1:0]) 
                    2'b00: begin 
                        wdata_o   <= {{16{mem_data_i[31]}}, mem_data_i[31:16]}; 
                        mem_sel_o <= 4'b1100; 
                    end 
                    2'b10: begin 
                        wdata_o   <= {{16{mem_data_i[15]}}, mem_data_i[15:0]}; 
                        mem_sel_o <= 4'b0011; 
                    end 
                    default: begin 
                        wdata_o   <= `ZeroWord; 
                    end 
                endcase 
            end
            `EXE_LHU_OP: begin            // lhu ָ�� 
                mem_addr_o <= mem_addr_i; 
                mem_we     <= `WriteDisable; 
                mem_ce_o   <= `ChipEnable; 
                case (mem_addr_i[1:0]) 
                    2'b00: begin 
                        wdata_o   <= {{16{1'b0}}, mem_data_i[31:16]}; 
                        mem_sel_o <= 4'b1100; 
                    end 
                    2'b10: begin 
                        wdata_o   <= {{16{1'b0}}, mem_data_i[15:0]}; 
                        mem_sel_o <= 4'b0011; 
                    end
                    default:       begin 
                        wdata_o   <= `ZeroWord; 
                    end 
                endcase 
            end
            `EXE_LW_OP: begin                   // lw ָ�� 
                mem_addr_o <= mem_addr_i; 
                mem_we     <= `WriteDisable; 
                wdata_o    <= mem_data_i; 
                mem_sel_o  <= 4'b1111; 
                mem_ce_o   <= `ChipEnable; 
            end 
            `EXE_LWL_OP: begin            // lwl ָ�� 
                mem_addr_o <= {mem_addr_i[31:2], 2'b00}; 
                mem_we     <= `WriteDisable; 
                mem_sel_o  <= 4'b1111; 
                mem_ce_o   <= `ChipEnable; 
                case (mem_addr_i[1:0]) 
                    2'b00: begin 
                        wdata_o <= mem_data_i[31:0]; 
                    end 
                    2'b01: begin 
                        wdata_o <= {mem_data_i[23:0], reg2_i[7:0]}; 
                    end 
                    2'b10: begin 
                        wdata_o <= {mem_data_i[15:0], reg2_i[15:0]}; 
                    end 
                    2'b11: begin 
                        wdata_o <= {mem_data_i[7:0], reg2_i[23:0]}; 
                    end 
                    default: begin 
                        wdata_o <= `ZeroWord; 
                    end 
                endcase 
            end
            `EXE_LWR_OP: begin             // lwr ָ�� 
                mem_addr_o <= {mem_addr_i[31:2], 2'b00}; 
                mem_we     <= `WriteDisable; 
                mem_sel_o  <= 4'b1111; 
                mem_ce_o   <= `ChipEnable; 
                case (mem_addr_i[1:0]) 
                    2'b00: begin 
                        wdata_o <= {reg2_i[31:8],mem_data_i[31:24]}; 
                    end
                    2'b01: begin 
                        wdata_o <= {reg2_i[31:16],mem_data_i[31:16]}; 
                    end 
                    2'b10: begin 
                        wdata_o <= {reg2_i[31:24],mem_data_i[31:8]}; 
                    end 
                    2'b11: begin 
                        wdata_o <= mem_data_i; 
                    end 
                    default: begin 
                        wdata_o <= `ZeroWord; 
                    end 
                endcase 
            end
            `EXE_LL_OP: begin               // ll ָ��ķô���� 
                mem_addr_o    <= mem_addr_i; 
                mem_we        <= `WriteDisable; 
                wdata_o       <= mem_data_i; 
                LLbit_we_o    <= 1'b1; 
                LLbit_value_o <= 1'b1; 
                mem_sel_o     <= 4'b1111; 
                mem_ce_o      <= `ChipEnable; 
            end
            `EXE_SB_OP: begin             // sb ָ�� 
                mem_addr_o <= mem_addr_i; 
                mem_we     <= `WriteEnable; 
                mem_data_o <= {reg2_i[7:0], reg2_i[7:0], reg2_i[7:0], reg2_i[7:0]}; 
                mem_ce_o   <= `ChipEnable; 
                case (mem_addr_i[1:0]) // ʵ���ϵ�ַֻ�и� 30 λ��Ч��Ϊ��� Wishbone ����
                    2'b00: begin 
                        mem_sel_o <= 4'b1000; 
                    end 
                    2'b01: begin 
                        mem_sel_o <= 4'b0100; 
                    end 
                    2'b10: begin 
                        mem_sel_o <= 4'b0010; 
                    end 
                    2'b11: begin 
                        mem_sel_o <= 4'b0001;  
                    end 
                    default: begin 
                        mem_sel_o <= 4'b0000; 
                    end 
                endcase 
            end
            `EXE_SH_OP: begin             // sh ָ�� 
                mem_addr_o <= mem_addr_i; 
                mem_we     <= `WriteEnable; 
                mem_data_o <= {reg2_i[15:0],reg2_i[15:0]}; 
                mem_ce_o   <= `ChipEnable; 
                case (mem_addr_i[1:0])
                    2'b00: begin 
                        mem_sel_o <= 4'b1100; 
                    end 
                    2'b10: begin 
                        mem_sel_o <= 4'b0011; 
                    end 
                    default: begin 
                        mem_sel_o <= 4'b0000; 
                    end 
                endcase 
            end
            `EXE_SW_OP: begin             // sw ָ�� 
                mem_addr_o <= mem_addr_i; 
                mem_we     <= `WriteEnable; 
                mem_data_o <= reg2_i; 
                mem_sel_o  <= 4'b1111; 
                mem_ce_o   <= `ChipEnable; 
            end
            `EXE_SWL_OP: begin             // swl ָ�� 
                mem_addr_o <= {mem_addr_i[31:2], 2'b00}; 
                mem_we     <= `WriteEnable; 
                mem_ce_o   <= `ChipEnable; 
                case (mem_addr_i[1:0]) 
                    2'b00: begin  
                        mem_sel_o <= 4'b1111; 
                        mem_data_o <= reg2_i; 
                    end 
                    2'b01: begin 
                        mem_sel_o <= 4'b0111; 
                        mem_data_o <= {zero32[7:0], reg2_i[31:8]}; 
                    end 
                    2'b10: begin 
                        mem_sel_o <= 4'b0011; 
                        mem_data_o <= {zero32[15:0], reg2_i[31:16]}; 
                    end 
                    2'b11: begin 
                        mem_sel_o <= 4'b0001; 
                        mem_data_o <= {zero32[23:0], reg2_i[31:24]}; 
                    end 
                    default: begin 
                        mem_sel_o <= 4'b0000; 
                    end 
                endcase 
            end
            `EXE_SWR_OP:  begin             // swr ָ�� 
                mem_addr_o <= {mem_addr_i[31:2], 2'b00}; 
                mem_we     <= `WriteEnable;
                mem_ce_o   <= `ChipEnable; 
                case (mem_addr_i[1:0]) 
                    2'b00: begin  
                        mem_sel_o  <= 4'b1000; 
                        mem_data_o <= {reg2_i[7:0], zero32[23:0]}; 
                    end 
                    2'b01: begin 
                        mem_sel_o  <= 4'b1100; 
                        mem_data_o <= {reg2_i[15:0],zero32[15:0]}; 
                    end 
                    2'b10: begin 
                        mem_sel_o  <= 4'b1110; 
                        mem_data_o <= {reg2_i[23:0],zero32[7:0]}; 
                    end 
                    2'b11: begin 
                        mem_sel_o  <= 4'b1111; 
                        mem_data_o <= reg2_i[31:0]; 
                    end 
                    default: begin 
                        mem_sel_o  <= 4'b0000; 
                    end 
                endcase 
            end
            `EXE_SC_OP: begin              // sc ָ��ķô���� 
                if(LLbit == 1'b1) begin 
                    LLbit_we_o    <= 1'b1; 
                    LLbit_value_o <= 1'b0; 
                    mem_addr_o    <= mem_addr_i; 
                    mem_we        <= `WriteEnable; 
                    mem_data_o    <= reg2_i; 
                    wdata_o       <= 32'b1; 
                    mem_sel_o     <= 4'b1111; 
                    mem_ce_o      <= `ChipEnable; 
                end 
                else begin 
                    wdata_o       <= 32'b0; 
                end 
            end
            default: begin 
                //do nothing 
            end
        endcase
    end     
end    

/**************************************************************** 
***********         ��һ�Σ��õ�CP0�мĴ���������ֵ        ********* 
*****************************************************************/

   // �õ� CP0 �� Status �Ĵ���������ֵ���������£� 
   // �жϵ�ǰ���ڻ�д�׶ε�ָ���Ƿ�Ҫд CP0 �� Status �Ĵ��������Ҫд����ôҪд 
   // ���ֵ���� Status �Ĵ���������ֵ����֮���� CP0 ģ��ͨ�� cp0_status_i �ӿ� 
   // ��������ݾ��� Status �Ĵ���������ֵ
   
always @ (*) begin 
    if(rst == `RstEnable) begin
        cp0_status <= `ZeroWord; 
    end 
    else if((wb_cp0_reg_we == `WriteEnable) && (wb_cp0_reg_write_addr == `CP0_REG_STATUS )) begin 
        cp0_status <= wb_cp0_reg_data; 
    end 
    else begin 
        cp0_status <= cp0_status_i; 
    end 
end

   // �õ� CP0 �� EPC �Ĵ���������ֵ���������£� 
   // �жϵ�ǰ���ڻ�д�׶ε�ָ���Ƿ�Ҫд CP0 �� EPC �Ĵ��������Ҫд����ôҪд�� 
   // ��ֵ���� EPC �Ĵ���������ֵ����֮���� CP0 ģ��ͨ�� cp0_epc_i �ӿڴ������ 
   // �ݾ��� EPC �Ĵ���������ֵ 
always @ (*) begin 
    if(rst == `RstEnable) begin 
        cp0_epc <= `ZeroWord; 
    end 
    else if((wb_cp0_reg_we == `WriteEnable) && (wb_cp0_reg_write_addr == `CP0_REG_EPC ))begin  
        cp0_epc <= wb_cp0_reg_data; 
    end 
    else begin 
        cp0_epc <= cp0_epc_i; 
    end 
end

    // �� EPC �Ĵ���������ֵͨ���ӿ� cp0_epc_o ��� 
    assign cp0_epc_o = cp0_epc;
   
   // �õ� CP0 �� Cause �Ĵ���������ֵ���������£� 
   // �жϵ�ǰ���ڻ�д�׶ε�ָ���Ƿ�Ҫд CP0 �� Cause �Ĵ��������Ҫд����ôҪд�� 
   // ��ֵ���� Cause �Ĵ���������ֵ������ע��һ�㣺Cause �Ĵ���ֻ�м����ֶ��ǿ�д 
   // �ġ���֮���� CP0 ģ��ͨ�� cp0_cause_i �ӿڴ�������ݾ��� Cause �Ĵ��������� 
   // ֵ 
always @ (*) begin 
    if(rst == `RstEnable) begin 
        cp0_cause <= `ZeroWord; 
    end 
    else if((wb_cp0_reg_we == `WriteEnable) && (wb_cp0_reg_write_addr == `CP0_REG_CAUSE )) begin 
        cp0_cause[9:8] <= wb_cp0_reg_data[9:8];  // IP[1:0] �ֶ��ǿ�д�� 
        cp0_cause[22]  <= wb_cp0_reg_data[22];   // WP �ֶ��ǿ�д�� 
        cp0_cause[23]  <= wb_cp0_reg_data[23];   // IV �ֶ��ǿ�д�� 
    end 
    else begin 
        cp0_cause      <= cp0_cause_i; 
    end 
end

/**************************************************************** 
***********           �ڶ��Σ��������յ��쳣����          ********* 
*****************************************************************/ 

always @ (*) begin 
    if(rst == `RstEnable) begin 
        excepttype_o <= `ZeroWord; 
    end 
    else begin 
        excepttype_o <= `ZeroWord; 
        if(current_inst_address_i != `ZeroWord) begin 
            if(((cp0_cause[15:8] & (cp0_status[15:8])) != 8'h00) && (cp0_status[1] == 1'b0) && (cp0_status[0] == 1'b1)) begin 
                excepttype_o <= 32'h00000001;            // interrupt 
            end 
            else if(excepttype_i[8]  == 1'b1) begin 
                excepttype_o <= 32'h00000008;            // syscall 
            end 
            else if(excepttype_i[9]  == 1'b1) begin 
                excepttype_o <= 32'h0000000a;            // inst_invalid 
            end 
            else if(excepttype_i[10] == 1'b1) begin 
                excepttype_o <= 32'h0000000d;            // trap 
            end 
            else if(excepttype_i[11] == 1'b1) begin   
                excepttype_o <= 32'h0000000c;            // ov 
            end 
            else if(excepttype_i[12] == 1'b1) begin   
                excepttype_o <= 32'h0000000e;            // eret 
            end 
            else if(excepttype_i[13] == 1'b1) begin
                excepttype_o <= 32'h00000009;            // break
            end
        end 
    end 
end

/**************************************************************** 
***********         �����Σ����������ݴ洢����д����        ********* 
*****************************************************************/ 
 
   // mem_we_o ��������ݴ洢������ʾ�Ƿ��Ƕ����ݴ洢����д������ 
   // ����������쳣����ô��Ҫȡ�������ݴ洢����д���� 
   assign mem_we_o = mem_we & (~(|excepttype_o));
   
   // һ�����ߴ���ÿһλ����������

endmodule
