`include "defines.vh"

module data_ram( 
       input  wire                   clk, 
       input  wire                   ce,        // ���ݴ洢��ʹ���ź�
       input  wire                   we,        // �Ƿ���д������Ϊ 1 ��ʾ��д����
       input  wire[`DataAddrBus]     addr,      // Ҫ���ʵĵ�ַ
       input  wire[3:0]              sel,       // �ֽ�ѡ���ź�
       input  wire[`DataBus]         data_i,    // Ҫд�������
       output reg [`DataBus]         data_o,    // ����������
       output [`DataBus]             seg7x16_data  // ������߶�����ܵ�����
);

       // �����ĸ��ֽ����� 
       reg[`ByteWidth]  data_mem0[0:`DataMemNum - 1]; 
       reg[`ByteWidth]  data_mem1[0:`DataMemNum - 1];
       reg[`ByteWidth]  data_mem2[0:`DataMemNum - 1]; 
       reg[`ByteWidth]  data_mem3[0:`DataMemNum - 1]; 
       
       // mem3 ��ʾģ 4 �� 0 �ĵ�ַ
       // mem2 ��ʾģ 4 �� 1 �ĵ�ַ
       // mem1 ��ʾģ 4 �� 2 �ĵ�ַ
       // mem0 ��ʾģ 4 �� 3 �ĵ�ַ
       
       assign seg7x16_data = {data_mem3[0], data_mem2[0], data_mem1[0], data_mem0[0]};
       
       // д���� 
        always @ (posedge clk) begin 
            if (ce == `ChipDisable) begin 
            // data_o <= ZeroWord; 
            end 
            else if(we == `WriteEnable) begin 
                if (sel[3] == 1'b1) begin // �ⲻ�����飡������������������ߵ�һλ�������� 3.2.1.0
                    data_mem3[addr[`DataMemNumLog2 + 1:2] - 17'b0_0100_0000_0000_0000] <= data_i[31:24]; // ���� 4 // �͵�ַ
                end 
                if (sel[2] == 1'b1) begin 
                    data_mem2[addr[`DataMemNumLog2 + 1:2] - 17'b0_0100_0000_0000_0000] <= data_i[23:16]; 
                end 
                if (sel[1] == 1'b1) begin 
                    data_mem1[addr[`DataMemNumLog2 + 1:2] - 17'b0_0100_0000_0000_0000] <= data_i[15:8]; 
                end 
                if (sel[0] == 1'b1) begin 
                    data_mem0[addr[`DataMemNumLog2 + 1:2] - 17'b0_0100_0000_0000_0000] <= data_i[7:0]; 
                end            
            end 
        end 
        
        // ������ ���� 0 1 2 3 ��ַ������
        always @ (*) begin 
            if (ce == `ChipDisable) begin 
                data_o <= `ZeroWord; 
            end 
            else if(we == `WriteDisable) begin // �� �� �� 0 1 2 3
                data_o <= {data_mem3[addr[`DataMemNumLog2 + 1:2] - 17'b0_0100_0000_0000_0000], 
                           data_mem2[addr[`DataMemNumLog2 + 1:2] - 17'b0_0100_0000_0000_0000], 
                           data_mem1[addr[`DataMemNumLog2 + 1:2] - 17'b0_0100_0000_0000_0000], 
                           data_mem0[addr[`DataMemNumLog2 + 1:2] - 17'b0_0100_0000_0000_0000]}; 
                           // - 17'b0_0100_0000_0000_0000 ����Ϊ MARS ���ݶ��Ǵ� 0x10010000 ��ʼ��
                           // 17'b0_0100_0000_0000_0000 �� 17'b1_0000_0000_0000_0000��0x10000�� ������λ������4���õ���
                           // �൱���� 19 λ��ַ���� 4 �õ� 17 λ��ַ���Ĵ�����ַ��������� 19 λ��ַ
                           // ���� MARS �е� 32 λ��ַ��32'b0001_0000_0000_0001_0000_0000_0000_0000��û��ȫ������
                           // ֻ���� 17'b1_0000_0000_0000_0000��0x10000��
            end 
            else begin 
                data_o <= `ZeroWord; 
            end 
        end

endmodule
