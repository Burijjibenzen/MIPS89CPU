`include "defines.vh"

module pc_reg( 
    input  wire              clk, 
    input  wire              rst, 
    input  wire[5:0]         stall, // ���Կ���ģ�� ctrl
    
    // ��������׶� ID ģ�����Ϣ 
    input wire               branch_flag_i, 
    input wire[`RegBus]      branch_target_address_i,
    
    input wire               flush,   // ��ˮ������ź�
    input wire[`RegBus]      new_pc,  // �쳣����������ڵ�ַ
    
    output reg[`InstAddrBus] pc, 
    output reg               ce   // ָ��洢��ʹ���ź�
);

always @ (posedge clk) begin 
    if (rst == `RstEnable) begin 
        ce <= `ChipDisable;       // ��λ��ʱ��ָ��洢������ 
    end 
    else begin
        ce <= `ChipEnable;        // ��λ������ָ��洢��ʹ�� 
    end 
end 

always @ (posedge clk) begin 
    if (ce == `ChipDisable) begin 
        pc <= 32'h30000000;       // ָ��洢�����õ�ʱ��PC Ϊ 0 
    end 
    else begin
        if (flush == 1'b1) begin
            // �����ź� flush Ϊ 1 ��ʾ�쳣���������� CTRL ģ��������쳣���� 
            // ������ڵ�ַ new_pc ��ȡִָ�� 
            pc <= new_pc;
        end
        else if (stall[0] == `NoStop) begin
            if (branch_flag_i == `Branch) begin 
                pc <= branch_target_address_i; 
            end
            else begin
                pc <= pc + 4'h4;
            end
        end
    end
end 

endmodule 