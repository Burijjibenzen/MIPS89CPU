`include "defines.vh"

module ctrl( 
    input wire          rst, 
    input wire          stallreq_from_id,   // ��������׶ε���ͣ���� 
    input wire          stallreq_from_ex,   // ����ִ�н׶ε���ͣ���� 
    
    // ���� MEM
    input wire[31:0]    excepttype_i,
    input wire[`RegBus] cp0_epc_i,
    
    output reg[`RegBus] new_pc,             // �쳣������ڵ�ַ 
    output reg          flush,              // �Ƿ������ˮ�� 
    
    output reg[5:0]     stall             
);

always @ (*) begin 
    if(rst == `RstEnable) begin 
        stall  <= 6'b000000; 
        flush  <= 1'b0; 
        new_pc <= `ZeroWord;
    end 
    else if(excepttype_i != `ZeroWord) begin  // ��Ϊ 0����ʾ�����쳣
        flush  <= 1'b1; 
        stall  <= 6'b000000;
        case (excepttype_i)
            32'h00000001: begin              // �ж� 
                new_pc <= 32'h00000020; 
            end
            32'h00000008: begin              // ϵͳ�����쳣 syscall 
                new_pc <= 32'h00400004;      // �ж����̵�ַ ��MARS��
            end
            32'h0000000a: begin              // ��Чָ���쳣 
                new_pc <= 32'h00400004; 
            end 
            32'h0000000d: begin              // �����쳣 
                new_pc <= 32'h00400004; 
            end 
            32'h0000000c: begin              // ����쳣 
                new_pc <= 32'h00400004; 
            end 
            32'h0000000e: begin              // �쳣����ָ�� eret 
                new_pc <= cp0_epc_i; 
            end 
            32'h00000009: begin              // �ϵ��쳣ָ�� break
                new_pc <= 32'h00400004;      // �Զ���
            end
            default: begin 
            end
        endcase
    end
    else if(stallreq_from_ex == `Stop) begin 
        stall <= 6'b001111; 
        flush <= 1'b0;
    end 
    else if(stallreq_from_id == `Stop) begin 
        stall <= 6'b000111; 
        flush <= 1'b0;
    end 
    else begin 
        stall  <= 6'b000000; 
        flush  <= 1'b0;
        new_pc <= `ZeroWord;
    end 
end

// stall[0] ��ʾȡָ��ַ PC �Ƿ񱣳ֲ��䣬Ϊ 1 ��ʾ���ֲ��䡣 
// stall[1] ��ʾ��ˮ��ȡָ�׶��Ƿ���ͣ��Ϊ 1 ��ʾ��ͣ�� 
// stall[2] ��ʾ��ˮ������׶��Ƿ���ͣ��Ϊ 1 ��ʾ��ͣ�� 
// stall[3] ��ʾ��ˮ��ִ�н׶��Ƿ���ͣ��Ϊ 1 ��ʾ��ͣ�� 
// stall[4] ��ʾ��ˮ�߷ô�׶��Ƿ���ͣ��Ϊ 1 ��ʾ��ͣ�� 
// stall[5] ��ʾ��ˮ�߻�д�׶��Ƿ���ͣ��Ϊ 1 ��ʾ��ͣ��

endmodule